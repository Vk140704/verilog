module and_gate(input i0,i1,output out);
 and g1(out,i0,i1);
 endmodule
