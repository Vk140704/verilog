module bufgate(input a,output y);
buf(y,a);
endmodule

