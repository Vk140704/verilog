// Code your testbench here
// or browse Examples
module lfsrtb;
reg clk,rst;
wire [3:0]op;
  lfsr lf1(.clk(clk),.rst(rst),.op(op));
  
  initial begin
    $dumpfile("lfsrtb.vcd");
    $dumpvars();
  end
  initial begin
    $monitor("op=%b",op);
    clk=0; rst=1;
    #5 rst=0;
    #50; $finish;
  end
  always #2 clk =~clk;
endmodule
