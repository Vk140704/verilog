module xorgate(input a,b,output out);
xor(out,a,b);
endmodule
