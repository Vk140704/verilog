module notgate(input a,output out);
not(out,a);
endmodule

