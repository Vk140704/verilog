module norgate (input a,b,output out);
nor(out,a,b);
endmodule
