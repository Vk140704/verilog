module ()
  
  endmodule
