module orgate(input a,b,output out);
or(out,a,b);
endmodule


