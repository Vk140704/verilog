module xnorgate(input a,b,output out);
xnor(out,a,b);
endmodule
