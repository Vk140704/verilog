module rcs(input[3:0] a,b,output [2:0]dif,output brw);
wire [2:0] b_out;

